//Verilog Code for AND Gate
module andgate(a,b,o);
 input a,b;
 output o;
  assign o=a&b;
endmodule
